
module ODDR(
    output wire Q,
    input wire D1, D2,
    input wire C,
    input wire CE, R,S
);

endmodule


module IBUFGDS (
    input wire I, IB,
    output wire O
);


endmodule
