
module system_wrapper
(
    inout wire [14:0]DDR_addr,
    inout wire [2:0]DDR_ba,
    inout wire DDR_cas_n,
    inout wire DDR_ck_n,
    inout wire DDR_ck_p,
    inout wire DDR_cke,
    inout wire DDR_cs_n,
    inout wire [3:0]DDR_dm,
    inout wire [31:0]DDR_dq,
    inout wire [3:0]DDR_dqs_n,
    inout wire [3:0]DDR_dqs_p,
    inout wire DDR_odt,
    inout wire DDR_ras_n,
    inout wire DDR_reset_n,
    inout wire DDR_we_n,
    inout wire FIXED_IO_ddr_vrn,
    inout wire FIXED_IO_ddr_vrp,
    inout wire [53:0]FIXED_IO_mio,
    inout wire FIXED_IO_ps_clk,
    inout wire FIXED_IO_ps_porb,
    inout wire FIXED_IO_ps_srstb,
    //axi signals
    output wire [31:0]M00_AXI_araddr,
    output wire [2:0]M00_AXI_arprot,
    input wire M00_AXI_arready,
    output wire M00_AXI_arvalid,
    output wire [31:0]M00_AXI_awaddr,
    output wire [2:0]M00_AXI_awprot,
    input wire M00_AXI_awready,
    output wire M00_AXI_awvalid,
    output wire M00_AXI_bready,
    input wire [1:0]M00_AXI_bresp,
    input wire M00_AXI_bvalid,
    input wire [31:0]M00_AXI_rdata,
    output wire M00_AXI_rready,
    input wire [1:0]M00_AXI_rresp,
    input wire M00_AXI_rvalid,
    output wire [31:0]M00_AXI_wdata,
    input wire M00_AXI_wready,
    output wire [3:0]M00_AXI_wstrb,
    output wire M00_AXI_wvalid,

    output wire [31:0]M01_AXI_araddr,
    output wire [2:0]M01_AXI_arprot,
    input wire M01_AXI_arready,
    output wire M01_AXI_arvalid,
    output wire [31:0]M01_AXI_awaddr,
    output wire [2:0]M01_AXI_awprot,
    input wire M01_AXI_awready,
    output wire M01_AXI_awvalid,
    output wire M01_AXI_bready,
    input wire [1:0]M01_AXI_bresp,
    input wire M01_AXI_bvalid,
    input wire [31:0]M01_AXI_rdata,
    output wire M01_AXI_rready,
    input wire [1:0]M01_AXI_rresp,
    input wire M01_AXI_rvalid,
    output wire [31:0]M01_AXI_wdata,
    input wire M01_AXI_wready,
    output wire [3:0]M01_AXI_wstrb,
    output wire M01_AXI_wvalid,

    output wire [31:0]M02_AXI_araddr,
    output wire [2:0]M02_AXI_arprot,
    input wire M02_AXI_arready,
    output wire M02_AXI_arvalid,
    output wire [31:0]M02_AXI_awaddr,
    output wire [2:0]M02_AXI_awprot,
    input wire M02_AXI_awready,
    output wire M02_AXI_awvalid,
    output wire M02_AXI_bready,
    input wire [1:0]M02_AXI_bresp,
    input wire M02_AXI_bvalid,
    input wire [31:0]M02_AXI_rdata,
    output wire M02_AXI_rready,
    input wire [1:0]M02_AXI_rresp,
    input wire M02_AXI_rvalid,
    output wire [31:0]M02_AXI_wdata,
    input wire M02_AXI_wready,
    output wire [3:0]M02_AXI_wstrb,
    output wire M02_AXI_wvalid,

    output wire [31:0]M03_AXI_araddr,
    output wire [2:0]M03_AXI_arprot,
    input wire M03_AXI_arready,
    output wire M03_AXI_arvalid,
    output wire [31:0]M03_AXI_awaddr,
    output wire [2:0]M03_AXI_awprot,
    input wire M03_AXI_awready,
    output wire M03_AXI_awvalid,
    output wire M03_AXI_bready,
    input wire [1:0]M03_AXI_bresp,
    input wire M03_AXI_bvalid,
    input wire [31:0]M03_AXI_rdata,
    output wire M03_AXI_rready,
    input wire [1:0]M03_AXI_rresp,
    input wire M03_AXI_rvalid,
    output wire [31:0]M03_AXI_wdata,
    input wire M03_AXI_wready,
    output wire [3:0]M03_AXI_wstrb,
    output wire M03_AXI_wvalid,
    
    output wire [31:0]M04_AXI_araddr,
    output wire [2:0]M04_AXI_arprot,
    input wire M04_AXI_arready,
    output wire M04_AXI_arvalid,
    output wire [31:0]M04_AXI_awaddr,
    output wire [2:0]M04_AXI_awprot,
    input wire M04_AXI_awready,
    output wire M04_AXI_awvalid,
    output wire M04_AXI_bready,
    input wire [1:0]M04_AXI_bresp,
    input wire M04_AXI_bvalid,
    input wire [31:0]M04_AXI_rdata,
    output wire M04_AXI_rready,
    input wire [1:0]M04_AXI_rresp,
    input wire M04_AXI_rvalid,
    output wire [31:0]M04_AXI_wdata,
    input wire M04_AXI_wready,
    output wire [3:0]M04_AXI_wstrb,
    output wire M04_AXI_wvalid,
    
    output wire [31:0]M05_AXI_araddr,
    output wire [2:0]M05_AXI_arprot,
    input wire M05_AXI_arready,
    output wire M05_AXI_arvalid,
    output wire [31:0]M05_AXI_awaddr,
    output wire [2:0]M05_AXI_awprot,
    input wire M05_AXI_awready,
    output wire M05_AXI_awvalid,
    output wire M05_AXI_bready,
    input wire [1:0]M05_AXI_bresp,
    input wire M05_AXI_bvalid,
    input wire [31:0]M05_AXI_rdata,
    output wire M05_AXI_rready,
    input wire [1:0]M05_AXI_rresp,
    input wire M05_AXI_rvalid,
    output wire [31:0]M05_AXI_wdata,
    input wire M05_AXI_wready,
    output wire [3:0]M05_AXI_wstrb,
    output wire M05_AXI_wvalid,
    
    output wire [31:0]M06_AXI_araddr,
    output wire [2:0]M06_AXI_arprot,
    input wire M06_AXI_arready,
    output wire M06_AXI_arvalid,
    output wire [31:0]M06_AXI_awaddr,
    output wire [2:0]M06_AXI_awprot,
    input wire M06_AXI_awready,
    output wire M06_AXI_awvalid,
    output wire M06_AXI_bready,
    input wire [1:0]M06_AXI_bresp,
    input wire M06_AXI_bvalid,
    input wire [31:0]M06_AXI_rdata,
    output wire M06_AXI_rready,
    input wire [1:0]M06_AXI_rresp,
    input wire M06_AXI_rvalid,
    output wire [31:0]M06_AXI_wdata,
    input wire M06_AXI_wready,
    output wire [3:0]M06_AXI_wstrb,
    output wire M06_AXI_wvalid,
    
    //clocks
    output wire adc_clk_out,
    output wire axi_clock
  );


endmodule
